module MicroCodeTableInner(input clk, input ce, input reset, input [7:0] IR, input [2:0] State, output reg [8:0] M);
  reg [8:0] L[0:2047];
  initial begin
L[0] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2] = 9'b00_10_10100; // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
L[3] = 9'b00_10_10100; // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
L[4] = 9'b00_10_10101; // P->[SP--]
L[5] = 9'b00_11_00011; // [VECT]->T
L[6] = 9'b10_11_10011; // [VECT]:T->PC
L[7] = 9'b00_00_00000; // []
L[8] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[9] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[10] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[11] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[12] = 9'b00_01_01011; // [A0]->AH,T->AL
L[13] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[14] = 9'b00_00_00000; // []
L[15] = 9'b00_00_00000; // []
L[16] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[17] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[18] = 9'b00_00_00000; // []
L[19] = 9'b00_00_00000; // []
L[20] = 9'b00_00_00000; // []
L[21] = 9'b00_00_00000; // []
L[22] = 9'b00_00_00000; // []
L[23] = 9'b00_00_00000; // []
L[24] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[25] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[26] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[27] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[28] = 9'b00_01_01011; // [A0]->AH,T->AL
L[29] = 9'b00_01_00011; // [A0]->T
L[30] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[31] = 9'b10_01_00101; // T->[A0]
L[32] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[33] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[34] = 9'b00_00_00000; // []
L[35] = 9'b00_00_00000; // []
L[36] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[37] = 9'b00_00_00000; // []
L[38] = 9'b00_00_00000; // []
L[39] = 9'b00_00_00000; // []
L[40] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[41] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[42] = 9'b00_00_00000; // []
L[43] = 9'b00_00_00000; // []
L[44] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[45] = 9'b00_00_00000; // []
L[46] = 9'b00_00_00000; // []
L[47] = 9'b00_00_00000; // []
L[48] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[49] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[50] = 9'b00_00_00000; // []
L[51] = 9'b00_00_00000; // []
L[52] = 9'b00_01_00011; // [A0]->T
L[53] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[54] = 9'b10_01_00101; // T->[A0]
L[55] = 9'b00_00_00000; // []
L[56] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[57] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[58] = 9'b00_00_00000; // []
L[59] = 9'b00_00_00000; // []
L[60] = 9'b00_01_00011; // [A0]->T
L[61] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[62] = 9'b10_01_00101; // T->[A0]
L[63] = 9'b00_00_00000; // []
L[64] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[65] = 9'b00_00_00011; // [PC]->
L[66] = 9'b10_10_01111; // P->[SP--]
L[67] = 9'b00_00_00000; // []
L[68] = 9'b00_00_00000; // []
L[69] = 9'b00_00_00000; // []
L[70] = 9'b00_00_00000; // []
L[71] = 9'b00_00_00000; // []
L[72] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[73] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[74] = 9'b00_00_00000; // []
L[75] = 9'b00_00_00000; // []
L[76] = 9'b00_00_00000; // []
L[77] = 9'b00_00_00000; // []
L[78] = 9'b00_00_00000; // []
L[79] = 9'b00_00_00000; // []
L[80] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[81] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[82] = 9'b00_00_00000; // []
L[83] = 9'b00_00_00000; // []
L[84] = 9'b00_00_00000; // []
L[85] = 9'b00_00_00000; // []
L[86] = 9'b00_00_00000; // []
L[87] = 9'b00_00_00000; // []
L[88] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[89] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[90] = 9'b00_00_00000; // []
L[91] = 9'b00_00_00000; // []
L[92] = 9'b00_00_00000; // []
L[93] = 9'b00_00_00000; // []
L[94] = 9'b00_00_00000; // []
L[95] = 9'b00_00_00000; // []
L[96] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[97] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[98] = 9'b11_00_00001; // [PC++]->AH
L[99] = 9'b00_00_00000; // []
L[100] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[101] = 9'b00_00_00000; // []
L[102] = 9'b00_00_00000; // []
L[103] = 9'b00_00_00000; // []
L[104] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[105] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[106] = 9'b11_00_00001; // [PC++]->AH
L[107] = 9'b00_00_00000; // []
L[108] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[109] = 9'b00_00_00000; // []
L[110] = 9'b00_00_00000; // []
L[111] = 9'b00_00_00000; // []
L[112] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[113] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[114] = 9'b11_00_00001; // [PC++]->AH
L[115] = 9'b00_00_00000; // []
L[116] = 9'b00_01_00011; // [A0]->T
L[117] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[118] = 9'b10_01_00101; // T->[A0]
L[119] = 9'b00_00_00000; // []
L[120] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[121] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[122] = 9'b11_00_00001; // [PC++]->AH
L[123] = 9'b00_00_00000; // []
L[124] = 9'b00_01_00011; // [A0]->T
L[125] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[126] = 9'b10_01_00101; // T->[A0]
L[127] = 9'b00_00_00000; // []
L[128] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[129] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[130] = 9'b11_00_10001; // PC+T->PC
L[131] = 9'b00_00_00000; // []
L[132] = 9'b10_00_00011; // ['NO-OP', '']
L[133] = 9'b00_00_00000; // []
L[134] = 9'b00_00_00000; // []
L[135] = 9'b00_00_00000; // []
L[136] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[137] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[138] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[139] = 9'b01_01_01100; // [A0]->AH,T+Y->AL
L[140] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[141] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[142] = 9'b00_00_00000; // []
L[143] = 9'b00_00_00000; // []
L[144] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[145] = 9'b10_00_00011; // ['NO-OP', '']
L[146] = 9'b00_00_00000; // []
L[147] = 9'b00_00_00000; // []
L[148] = 9'b00_00_00000; // []
L[149] = 9'b00_00_00000; // []
L[150] = 9'b00_00_00000; // []
L[151] = 9'b00_00_00000; // []
L[152] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[153] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[154] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[155] = 9'b00_01_01100; // [A0]->AH,T+Y->AL
L[156] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[157] = 9'b00_01_00011; // [A0]->T
L[158] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[159] = 9'b10_01_00101; // T->[A0]
L[160] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[161] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[162] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[163] = 9'b00_00_00000; // []
L[164] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[165] = 9'b00_00_00000; // []
L[166] = 9'b00_00_00000; // []
L[167] = 9'b00_00_00000; // []
L[168] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[169] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[170] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[171] = 9'b00_00_00000; // []
L[172] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[173] = 9'b00_00_00000; // []
L[174] = 9'b00_00_00000; // []
L[175] = 9'b00_00_00000; // []
L[176] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[177] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[178] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[179] = 9'b00_00_00000; // []
L[180] = 9'b00_01_00011; // [A0]->T
L[181] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[182] = 9'b10_01_00101; // T->[A0]
L[183] = 9'b00_00_00000; // []
L[184] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[185] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[186] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[187] = 9'b00_00_00000; // []
L[188] = 9'b00_01_00011; // [A0]->T
L[189] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[190] = 9'b10_01_00101; // T->[A0]
L[191] = 9'b00_00_00000; // []
L[192] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[193] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[194] = 9'b00_00_00000; // []
L[195] = 9'b00_00_00000; // []
L[196] = 9'b00_00_00000; // []
L[197] = 9'b00_00_00000; // []
L[198] = 9'b00_00_00000; // []
L[199] = 9'b00_00_00000; // []
L[200] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[201] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[202] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[203] = 9'b00_00_00000; // []
L[204] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[205] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[206] = 9'b00_00_00000; // []
L[207] = 9'b00_00_00000; // []
L[208] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[209] = 9'b10_00_00011; // ['NO-OP', '']
L[210] = 9'b00_00_00000; // []
L[211] = 9'b00_00_00000; // []
L[212] = 9'b00_00_00000; // []
L[213] = 9'b00_00_00000; // []
L[214] = 9'b00_00_00000; // []
L[215] = 9'b00_00_00000; // []
L[216] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[217] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[218] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[219] = 9'b00_00_00000; // []
L[220] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[221] = 9'b00_01_00011; // [A0]->T
L[222] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[223] = 9'b10_01_00101; // T->[A0]
L[224] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[225] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[226] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[227] = 9'b00_00_00000; // []
L[228] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[229] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[230] = 9'b00_00_00000; // []
L[231] = 9'b00_00_00000; // []
L[232] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[233] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[234] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[235] = 9'b00_00_00000; // []
L[236] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[237] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[238] = 9'b00_00_00000; // []
L[239] = 9'b00_00_00000; // []
L[240] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[241] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[242] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[243] = 9'b00_00_00000; // []
L[244] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[245] = 9'b00_01_00011; // [A0]->T
L[246] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[247] = 9'b10_01_00101; // T->[A0]
L[248] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[249] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[250] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[251] = 9'b00_00_00000; // []
L[252] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[253] = 9'b00_01_00011; // [A0]->T
L[254] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[255] = 9'b10_01_00101; // T->[A0]
L[256] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[257] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[258] = 9'b00_10_10100; // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
L[259] = 9'b00_10_10100; // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
L[260] = 9'b00_10_00111; // KEEP_AC
L[261] = 9'b10_00_10011; // [PC]:T->PC
L[262] = 9'b00_00_00000; // []
L[263] = 9'b00_00_00000; // []
L[264] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[265] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[266] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[267] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[268] = 9'b00_01_01011; // [A0]->AH,T->AL
L[269] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[270] = 9'b00_00_00000; // []
L[271] = 9'b00_00_00000; // []
L[272] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[273] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[274] = 9'b00_00_00000; // []
L[275] = 9'b00_00_00000; // []
L[276] = 9'b00_00_00000; // []
L[277] = 9'b00_00_00000; // []
L[278] = 9'b00_00_00000; // []
L[279] = 9'b00_00_00000; // []
L[280] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[281] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[282] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[283] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[284] = 9'b00_01_01011; // [A0]->AH,T->AL
L[285] = 9'b00_01_00011; // [A0]->T
L[286] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[287] = 9'b10_01_00101; // T->[A0]
L[288] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[289] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[290] = 9'b00_00_00000; // []
L[291] = 9'b00_00_00000; // []
L[292] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[293] = 9'b00_00_00000; // []
L[294] = 9'b00_00_00000; // []
L[295] = 9'b00_00_00000; // []
L[296] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[297] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[298] = 9'b00_00_00000; // []
L[299] = 9'b00_00_00000; // []
L[300] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[301] = 9'b00_00_00000; // []
L[302] = 9'b00_00_00000; // []
L[303] = 9'b00_00_00000; // []
L[304] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[305] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[306] = 9'b00_00_00000; // []
L[307] = 9'b00_00_00000; // []
L[308] = 9'b00_01_00011; // [A0]->T
L[309] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[310] = 9'b10_01_00101; // T->[A0]
L[311] = 9'b00_00_00000; // []
L[312] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[313] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[314] = 9'b00_00_00000; // []
L[315] = 9'b00_00_00000; // []
L[316] = 9'b00_01_00011; // [A0]->T
L[317] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[318] = 9'b10_01_00101; // T->[A0]
L[319] = 9'b00_00_00000; // []
L[320] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[321] = 9'b00_00_00011; // [PC]->
L[322] = 9'b00_10_10000; // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
L[323] = 9'b10_10_00010; // ['ALU([SP])->A', '[SP]->P']
L[324] = 9'b00_00_00000; // []
L[325] = 9'b00_00_00000; // []
L[326] = 9'b00_00_00000; // []
L[327] = 9'b00_00_00000; // []
L[328] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[329] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[330] = 9'b00_00_00000; // []
L[331] = 9'b00_00_00000; // []
L[332] = 9'b00_00_00000; // []
L[333] = 9'b00_00_00000; // []
L[334] = 9'b00_00_00000; // []
L[335] = 9'b00_00_00000; // []
L[336] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[337] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[338] = 9'b00_00_00000; // []
L[339] = 9'b00_00_00000; // []
L[340] = 9'b00_00_00000; // []
L[341] = 9'b00_00_00000; // []
L[342] = 9'b00_00_00000; // []
L[343] = 9'b00_00_00000; // []
L[344] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[345] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[346] = 9'b00_00_00000; // []
L[347] = 9'b00_00_00000; // []
L[348] = 9'b00_00_00000; // []
L[349] = 9'b00_00_00000; // []
L[350] = 9'b00_00_00000; // []
L[351] = 9'b00_00_00000; // []
L[352] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[353] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[354] = 9'b11_00_00001; // [PC++]->AH
L[355] = 9'b00_00_00000; // []
L[356] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[357] = 9'b00_00_00000; // []
L[358] = 9'b00_00_00000; // []
L[359] = 9'b00_00_00000; // []
L[360] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[361] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[362] = 9'b11_00_00001; // [PC++]->AH
L[363] = 9'b00_00_00000; // []
L[364] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[365] = 9'b00_00_00000; // []
L[366] = 9'b00_00_00000; // []
L[367] = 9'b00_00_00000; // []
L[368] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[369] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[370] = 9'b11_00_00001; // [PC++]->AH
L[371] = 9'b00_00_00000; // []
L[372] = 9'b00_01_00011; // [A0]->T
L[373] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[374] = 9'b10_01_00101; // T->[A0]
L[375] = 9'b00_00_00000; // []
L[376] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[377] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[378] = 9'b11_00_00001; // [PC++]->AH
L[379] = 9'b00_00_00000; // []
L[380] = 9'b00_01_00011; // [A0]->T
L[381] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[382] = 9'b10_01_00101; // T->[A0]
L[383] = 9'b00_00_00000; // []
L[384] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[385] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[386] = 9'b11_00_10001; // PC+T->PC
L[387] = 9'b00_00_00000; // []
L[388] = 9'b10_00_00011; // ['NO-OP', '']
L[389] = 9'b00_00_00000; // []
L[390] = 9'b00_00_00000; // []
L[391] = 9'b00_00_00000; // []
L[392] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[393] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[394] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[395] = 9'b01_01_01100; // [A0]->AH,T+Y->AL
L[396] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[397] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[398] = 9'b00_00_00000; // []
L[399] = 9'b00_00_00000; // []
L[400] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[401] = 9'b10_00_00011; // ['NO-OP', '']
L[402] = 9'b00_00_00000; // []
L[403] = 9'b00_00_00000; // []
L[404] = 9'b00_00_00000; // []
L[405] = 9'b00_00_00000; // []
L[406] = 9'b00_00_00000; // []
L[407] = 9'b00_00_00000; // []
L[408] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[409] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[410] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[411] = 9'b00_01_01100; // [A0]->AH,T+Y->AL
L[412] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[413] = 9'b00_01_00011; // [A0]->T
L[414] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[415] = 9'b10_01_00101; // T->[A0]
L[416] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[417] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[418] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[419] = 9'b00_00_00000; // []
L[420] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[421] = 9'b00_00_00000; // []
L[422] = 9'b00_00_00000; // []
L[423] = 9'b00_00_00000; // []
L[424] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[425] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[426] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[427] = 9'b00_00_00000; // []
L[428] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[429] = 9'b00_00_00000; // []
L[430] = 9'b00_00_00000; // []
L[431] = 9'b00_00_00000; // []
L[432] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[433] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[434] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[435] = 9'b00_00_00000; // []
L[436] = 9'b00_01_00011; // [A0]->T
L[437] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[438] = 9'b10_01_00101; // T->[A0]
L[439] = 9'b00_00_00000; // []
L[440] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[441] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[442] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[443] = 9'b00_00_00000; // []
L[444] = 9'b00_01_00011; // [A0]->T
L[445] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[446] = 9'b10_01_00101; // T->[A0]
L[447] = 9'b00_00_00000; // []
L[448] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[449] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[450] = 9'b00_00_00000; // []
L[451] = 9'b00_00_00000; // []
L[452] = 9'b00_00_00000; // []
L[453] = 9'b00_00_00000; // []
L[454] = 9'b00_00_00000; // []
L[455] = 9'b00_00_00000; // []
L[456] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[457] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[458] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[459] = 9'b00_00_00000; // []
L[460] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[461] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[462] = 9'b00_00_00000; // []
L[463] = 9'b00_00_00000; // []
L[464] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[465] = 9'b10_00_00011; // ['NO-OP', '']
L[466] = 9'b00_00_00000; // []
L[467] = 9'b00_00_00000; // []
L[468] = 9'b00_00_00000; // []
L[469] = 9'b00_00_00000; // []
L[470] = 9'b00_00_00000; // []
L[471] = 9'b00_00_00000; // []
L[472] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[473] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[474] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[475] = 9'b00_00_00000; // []
L[476] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[477] = 9'b00_01_00011; // [A0]->T
L[478] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[479] = 9'b10_01_00101; // T->[A0]
L[480] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[481] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[482] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[483] = 9'b00_00_00000; // []
L[484] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[485] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[486] = 9'b00_00_00000; // []
L[487] = 9'b00_00_00000; // []
L[488] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[489] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[490] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[491] = 9'b00_00_00000; // []
L[492] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[493] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[494] = 9'b00_00_00000; // []
L[495] = 9'b00_00_00000; // []
L[496] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[497] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[498] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[499] = 9'b00_00_00000; // []
L[500] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[501] = 9'b00_01_00011; // [A0]->T
L[502] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[503] = 9'b10_01_00101; // T->[A0]
L[504] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[505] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[506] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[507] = 9'b00_00_00000; // []
L[508] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[509] = 9'b00_01_00011; // [A0]->T
L[510] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[511] = 9'b10_01_00101; // T->[A0]
L[512] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[513] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[514] = 9'b00_10_10000; // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
L[515] = 9'b00_10_10110; // [SP]->P,SP+1->SP
L[516] = 9'b00_10_10000; // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
L[517] = 9'b10_10_10011; // [SP]:T->PC
L[518] = 9'b00_00_00000; // []
L[519] = 9'b00_00_00000; // []
L[520] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[521] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[522] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[523] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[524] = 9'b00_01_01011; // [A0]->AH,T->AL
L[525] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[526] = 9'b00_00_00000; // []
L[527] = 9'b00_00_00000; // []
L[528] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[529] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[530] = 9'b00_00_00000; // []
L[531] = 9'b00_00_00000; // []
L[532] = 9'b00_00_00000; // []
L[533] = 9'b00_00_00000; // []
L[534] = 9'b00_00_00000; // []
L[535] = 9'b00_00_00000; // []
L[536] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[537] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[538] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[539] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[540] = 9'b00_01_01011; // [A0]->AH,T->AL
L[541] = 9'b00_01_00011; // [A0]->T
L[542] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[543] = 9'b10_01_00101; // T->[A0]
L[544] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[545] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[546] = 9'b00_00_00000; // []
L[547] = 9'b00_00_00000; // []
L[548] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[549] = 9'b00_00_00000; // []
L[550] = 9'b00_00_00000; // []
L[551] = 9'b00_00_00000; // []
L[552] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[553] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[554] = 9'b00_00_00000; // []
L[555] = 9'b00_00_00000; // []
L[556] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[557] = 9'b00_00_00000; // []
L[558] = 9'b00_00_00000; // []
L[559] = 9'b00_00_00000; // []
L[560] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[561] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[562] = 9'b00_00_00000; // []
L[563] = 9'b00_00_00000; // []
L[564] = 9'b00_01_00011; // [A0]->T
L[565] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[566] = 9'b10_01_00101; // T->[A0]
L[567] = 9'b00_00_00000; // []
L[568] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[569] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[570] = 9'b00_00_00000; // []
L[571] = 9'b00_00_00000; // []
L[572] = 9'b00_01_00011; // [A0]->T
L[573] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[574] = 9'b10_01_00101; // T->[A0]
L[575] = 9'b00_00_00000; // []
L[576] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[577] = 9'b00_00_00011; // [PC]->
L[578] = 9'b10_10_01110; // ALU(A)->[SP--]
L[579] = 9'b00_00_00000; // []
L[580] = 9'b00_00_00000; // []
L[581] = 9'b00_00_00000; // []
L[582] = 9'b00_00_00000; // []
L[583] = 9'b00_00_00000; // []
L[584] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[585] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[586] = 9'b00_00_00000; // []
L[587] = 9'b00_00_00000; // []
L[588] = 9'b00_00_00000; // []
L[589] = 9'b00_00_00000; // []
L[590] = 9'b00_00_00000; // []
L[591] = 9'b00_00_00000; // []
L[592] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[593] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[594] = 9'b00_00_00000; // []
L[595] = 9'b00_00_00000; // []
L[596] = 9'b00_00_00000; // []
L[597] = 9'b00_00_00000; // []
L[598] = 9'b00_00_00000; // []
L[599] = 9'b00_00_00000; // []
L[600] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[601] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[602] = 9'b00_00_00000; // []
L[603] = 9'b00_00_00000; // []
L[604] = 9'b00_00_00000; // []
L[605] = 9'b00_00_00000; // []
L[606] = 9'b00_00_00000; // []
L[607] = 9'b00_00_00000; // []
L[608] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[609] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[610] = 9'b00_00_00000; // []
L[611] = 9'b00_00_00000; // []
L[612] = 9'b10_00_10011; // [PC]:T->PC
L[613] = 9'b00_00_00000; // []
L[614] = 9'b00_00_00000; // []
L[615] = 9'b00_00_00000; // []
L[616] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[617] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[618] = 9'b11_00_00001; // [PC++]->AH
L[619] = 9'b00_00_00000; // []
L[620] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[621] = 9'b00_00_00000; // []
L[622] = 9'b00_00_00000; // []
L[623] = 9'b00_00_00000; // []
L[624] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[625] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[626] = 9'b11_00_00001; // [PC++]->AH
L[627] = 9'b00_00_00000; // []
L[628] = 9'b00_01_00011; // [A0]->T
L[629] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[630] = 9'b10_01_00101; // T->[A0]
L[631] = 9'b00_00_00000; // []
L[632] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[633] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[634] = 9'b11_00_00001; // [PC++]->AH
L[635] = 9'b00_00_00000; // []
L[636] = 9'b00_01_00011; // [A0]->T
L[637] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[638] = 9'b10_01_00101; // T->[A0]
L[639] = 9'b00_00_00000; // []
L[640] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[641] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[642] = 9'b11_00_10001; // PC+T->PC
L[643] = 9'b00_00_00000; // []
L[644] = 9'b10_00_00011; // ['NO-OP', '']
L[645] = 9'b00_00_00000; // []
L[646] = 9'b00_00_00000; // []
L[647] = 9'b00_00_00000; // []
L[648] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[649] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[650] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[651] = 9'b01_01_01100; // [A0]->AH,T+Y->AL
L[652] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[653] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[654] = 9'b00_00_00000; // []
L[655] = 9'b00_00_00000; // []
L[656] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[657] = 9'b10_00_00011; // ['NO-OP', '']
L[658] = 9'b00_00_00000; // []
L[659] = 9'b00_00_00000; // []
L[660] = 9'b00_00_00000; // []
L[661] = 9'b00_00_00000; // []
L[662] = 9'b00_00_00000; // []
L[663] = 9'b00_00_00000; // []
L[664] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[665] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[666] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[667] = 9'b00_01_01100; // [A0]->AH,T+Y->AL
L[668] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[669] = 9'b00_01_00011; // [A0]->T
L[670] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[671] = 9'b10_01_00101; // T->[A0]
L[672] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[673] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[674] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[675] = 9'b00_00_00000; // []
L[676] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[677] = 9'b00_00_00000; // []
L[678] = 9'b00_00_00000; // []
L[679] = 9'b00_00_00000; // []
L[680] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[681] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[682] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[683] = 9'b00_00_00000; // []
L[684] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[685] = 9'b00_00_00000; // []
L[686] = 9'b00_00_00000; // []
L[687] = 9'b00_00_00000; // []
L[688] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[689] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[690] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[691] = 9'b00_00_00000; // []
L[692] = 9'b00_01_00011; // [A0]->T
L[693] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[694] = 9'b10_01_00101; // T->[A0]
L[695] = 9'b00_00_00000; // []
L[696] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[697] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[698] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[699] = 9'b00_00_00000; // []
L[700] = 9'b00_01_00011; // [A0]->T
L[701] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[702] = 9'b10_01_00101; // T->[A0]
L[703] = 9'b00_00_00000; // []
L[704] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[705] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[706] = 9'b00_00_00000; // []
L[707] = 9'b00_00_00000; // []
L[708] = 9'b00_00_00000; // []
L[709] = 9'b00_00_00000; // []
L[710] = 9'b00_00_00000; // []
L[711] = 9'b00_00_00000; // []
L[712] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[713] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[714] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[715] = 9'b00_00_00000; // []
L[716] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[717] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[718] = 9'b00_00_00000; // []
L[719] = 9'b00_00_00000; // []
L[720] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[721] = 9'b10_00_00011; // ['NO-OP', '']
L[722] = 9'b00_00_00000; // []
L[723] = 9'b00_00_00000; // []
L[724] = 9'b00_00_00000; // []
L[725] = 9'b00_00_00000; // []
L[726] = 9'b00_00_00000; // []
L[727] = 9'b00_00_00000; // []
L[728] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[729] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[730] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[731] = 9'b00_00_00000; // []
L[732] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[733] = 9'b00_01_00011; // [A0]->T
L[734] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[735] = 9'b10_01_00101; // T->[A0]
L[736] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[737] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[738] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[739] = 9'b00_00_00000; // []
L[740] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[741] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[742] = 9'b00_00_00000; // []
L[743] = 9'b00_00_00000; // []
L[744] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[745] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[746] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[747] = 9'b00_00_00000; // []
L[748] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[749] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[750] = 9'b00_00_00000; // []
L[751] = 9'b00_00_00000; // []
L[752] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[753] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[754] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[755] = 9'b00_00_00000; // []
L[756] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[757] = 9'b00_01_00011; // [A0]->T
L[758] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[759] = 9'b10_01_00101; // T->[A0]
L[760] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[761] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[762] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[763] = 9'b00_00_00000; // []
L[764] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[765] = 9'b00_01_00011; // [A0]->T
L[766] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[767] = 9'b10_01_00101; // T->[A0]
L[768] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[769] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[770] = 9'b11_10_10000; // SP+1->SP
L[771] = 9'b00_00_00000; // []
L[772] = 9'b00_10_10000; // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
L[773] = 9'b00_10_10011; // [SP]:T->PC
L[774] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[775] = 9'b00_00_00000; // []
L[776] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[777] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[778] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[779] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[780] = 9'b00_01_01011; // [A0]->AH,T->AL
L[781] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[782] = 9'b00_00_00000; // []
L[783] = 9'b00_00_00000; // []
L[784] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[785] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[786] = 9'b00_00_00000; // []
L[787] = 9'b00_00_00000; // []
L[788] = 9'b00_00_00000; // []
L[789] = 9'b00_00_00000; // []
L[790] = 9'b00_00_00000; // []
L[791] = 9'b00_00_00000; // []
L[792] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[793] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[794] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[795] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[796] = 9'b00_01_01011; // [A0]->AH,T->AL
L[797] = 9'b00_01_00011; // [A0]->T
L[798] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[799] = 9'b10_01_00101; // T->[A0]
L[800] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[801] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[802] = 9'b00_00_00000; // []
L[803] = 9'b00_00_00000; // []
L[804] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[805] = 9'b00_00_00000; // []
L[806] = 9'b00_00_00000; // []
L[807] = 9'b00_00_00000; // []
L[808] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[809] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[810] = 9'b00_00_00000; // []
L[811] = 9'b00_00_00000; // []
L[812] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[813] = 9'b00_00_00000; // []
L[814] = 9'b00_00_00000; // []
L[815] = 9'b00_00_00000; // []
L[816] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[817] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[818] = 9'b00_00_00000; // []
L[819] = 9'b00_00_00000; // []
L[820] = 9'b00_01_00011; // [A0]->T
L[821] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[822] = 9'b10_01_00101; // T->[A0]
L[823] = 9'b00_00_00000; // []
L[824] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[825] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[826] = 9'b00_00_00000; // []
L[827] = 9'b00_00_00000; // []
L[828] = 9'b00_01_00011; // [A0]->T
L[829] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[830] = 9'b10_01_00101; // T->[A0]
L[831] = 9'b00_00_00000; // []
L[832] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[833] = 9'b00_00_00011; // [PC]->
L[834] = 9'b00_10_10000; // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
L[835] = 9'b10_10_00010; // ['ALU([SP])->A', '[SP]->P']
L[836] = 9'b00_00_00000; // []
L[837] = 9'b00_00_00000; // []
L[838] = 9'b00_00_00000; // []
L[839] = 9'b00_00_00000; // []
L[840] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[841] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[842] = 9'b00_00_00000; // []
L[843] = 9'b00_00_00000; // []
L[844] = 9'b00_00_00000; // []
L[845] = 9'b00_00_00000; // []
L[846] = 9'b00_00_00000; // []
L[847] = 9'b00_00_00000; // []
L[848] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[849] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[850] = 9'b00_00_00000; // []
L[851] = 9'b00_00_00000; // []
L[852] = 9'b00_00_00000; // []
L[853] = 9'b00_00_00000; // []
L[854] = 9'b00_00_00000; // []
L[855] = 9'b00_00_00000; // []
L[856] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[857] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[858] = 9'b00_00_00000; // []
L[859] = 9'b00_00_00000; // []
L[860] = 9'b00_00_00000; // []
L[861] = 9'b00_00_00000; // []
L[862] = 9'b00_00_00000; // []
L[863] = 9'b00_00_00000; // []
L[864] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[865] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[866] = 9'b00_00_00001; // [PC++]->AH
L[867] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[868] = 9'b10_01_10011; // [A0]:T->PC
L[869] = 9'b00_00_00000; // []
L[870] = 9'b00_00_00000; // []
L[871] = 9'b00_00_00000; // []
L[872] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[873] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[874] = 9'b11_00_00001; // [PC++]->AH
L[875] = 9'b00_00_00000; // []
L[876] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[877] = 9'b00_00_00000; // []
L[878] = 9'b00_00_00000; // []
L[879] = 9'b00_00_00000; // []
L[880] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[881] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[882] = 9'b11_00_00001; // [PC++]->AH
L[883] = 9'b00_00_00000; // []
L[884] = 9'b00_01_00011; // [A0]->T
L[885] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[886] = 9'b10_01_00101; // T->[A0]
L[887] = 9'b00_00_00000; // []
L[888] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[889] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[890] = 9'b11_00_00001; // [PC++]->AH
L[891] = 9'b00_00_00000; // []
L[892] = 9'b00_01_00011; // [A0]->T
L[893] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[894] = 9'b10_01_00101; // T->[A0]
L[895] = 9'b00_00_00000; // []
L[896] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[897] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[898] = 9'b11_00_10001; // PC+T->PC
L[899] = 9'b00_00_00000; // []
L[900] = 9'b10_00_00011; // ['NO-OP', '']
L[901] = 9'b00_00_00000; // []
L[902] = 9'b00_00_00000; // []
L[903] = 9'b00_00_00000; // []
L[904] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[905] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[906] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[907] = 9'b01_01_01100; // [A0]->AH,T+Y->AL
L[908] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[909] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[910] = 9'b00_00_00000; // []
L[911] = 9'b00_00_00000; // []
L[912] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[913] = 9'b10_00_00011; // ['NO-OP', '']
L[914] = 9'b00_00_00000; // []
L[915] = 9'b00_00_00000; // []
L[916] = 9'b00_00_00000; // []
L[917] = 9'b00_00_00000; // []
L[918] = 9'b00_00_00000; // []
L[919] = 9'b00_00_00000; // []
L[920] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[921] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[922] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[923] = 9'b00_01_01100; // [A0]->AH,T+Y->AL
L[924] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[925] = 9'b00_01_00011; // [A0]->T
L[926] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[927] = 9'b10_01_00101; // T->[A0]
L[928] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[929] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[930] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[931] = 9'b00_00_00000; // []
L[932] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[933] = 9'b00_00_00000; // []
L[934] = 9'b00_00_00000; // []
L[935] = 9'b00_00_00000; // []
L[936] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[937] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[938] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[939] = 9'b00_00_00000; // []
L[940] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[941] = 9'b00_00_00000; // []
L[942] = 9'b00_00_00000; // []
L[943] = 9'b00_00_00000; // []
L[944] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[945] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[946] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[947] = 9'b00_00_00000; // []
L[948] = 9'b00_01_00011; // [A0]->T
L[949] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[950] = 9'b10_01_00101; // T->[A0]
L[951] = 9'b00_00_00000; // []
L[952] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[953] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[954] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[955] = 9'b00_00_00000; // []
L[956] = 9'b00_01_00011; // [A0]->T
L[957] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[958] = 9'b10_01_00101; // T->[A0]
L[959] = 9'b00_00_00000; // []
L[960] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[961] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[962] = 9'b00_00_00000; // []
L[963] = 9'b00_00_00000; // []
L[964] = 9'b00_00_00000; // []
L[965] = 9'b00_00_00000; // []
L[966] = 9'b00_00_00000; // []
L[967] = 9'b00_00_00000; // []
L[968] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[969] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[970] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[971] = 9'b00_00_00000; // []
L[972] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[973] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[974] = 9'b00_00_00000; // []
L[975] = 9'b00_00_00000; // []
L[976] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[977] = 9'b10_00_00011; // ['NO-OP', '']
L[978] = 9'b00_00_00000; // []
L[979] = 9'b00_00_00000; // []
L[980] = 9'b00_00_00000; // []
L[981] = 9'b00_00_00000; // []
L[982] = 9'b00_00_00000; // []
L[983] = 9'b00_00_00000; // []
L[984] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[985] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[986] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[987] = 9'b00_00_00000; // []
L[988] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[989] = 9'b00_01_00011; // [A0]->T
L[990] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[991] = 9'b10_01_00101; // T->[A0]
L[992] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[993] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[994] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[995] = 9'b00_00_00000; // []
L[996] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[997] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[998] = 9'b00_00_00000; // []
L[999] = 9'b00_00_00000; // []
L[1000] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1001] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1002] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1003] = 9'b00_00_00000; // []
L[1004] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1005] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1006] = 9'b00_00_00000; // []
L[1007] = 9'b00_00_00000; // []
L[1008] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1009] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1010] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1011] = 9'b00_00_00000; // []
L[1012] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1013] = 9'b00_01_00011; // [A0]->T
L[1014] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1015] = 9'b10_01_00101; // T->[A0]
L[1016] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1017] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1018] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1019] = 9'b00_00_00000; // []
L[1020] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1021] = 9'b00_01_00011; // [A0]->T
L[1022] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1023] = 9'b10_01_00101; // T->[A0]
L[1024] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1025] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1026] = 9'b00_00_00000; // []
L[1027] = 9'b00_00_00000; // []
L[1028] = 9'b00_00_00000; // []
L[1029] = 9'b00_00_00000; // []
L[1030] = 9'b00_00_00000; // []
L[1031] = 9'b00_00_00000; // []
L[1032] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1033] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1034] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[1035] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1036] = 9'b00_01_01011; // [A0]->AH,T->AL
L[1037] = 9'b10_01_00110; // ALU()->[A0]
L[1038] = 9'b00_00_00000; // []
L[1039] = 9'b00_00_00000; // []
L[1040] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1041] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1042] = 9'b00_00_00000; // []
L[1043] = 9'b00_00_00000; // []
L[1044] = 9'b00_00_00000; // []
L[1045] = 9'b00_00_00000; // []
L[1046] = 9'b00_00_00000; // []
L[1047] = 9'b00_00_00000; // []
L[1048] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1049] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1050] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[1051] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1052] = 9'b00_01_01011; // [A0]->AH,T->AL
L[1053] = 9'b10_01_00110; // ALU()->[A0]
L[1054] = 9'b00_00_00000; // []
L[1055] = 9'b00_00_00000; // []
L[1056] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1057] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1058] = 9'b00_00_00000; // []
L[1059] = 9'b00_00_00000; // []
L[1060] = 9'b10_01_00110; // ALU()->[A0]
L[1061] = 9'b00_00_00000; // []
L[1062] = 9'b00_00_00000; // []
L[1063] = 9'b00_00_00000; // []
L[1064] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1065] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1066] = 9'b00_00_00000; // []
L[1067] = 9'b00_00_00000; // []
L[1068] = 9'b10_01_00110; // ALU()->[A0]
L[1069] = 9'b00_00_00000; // []
L[1070] = 9'b00_00_00000; // []
L[1071] = 9'b00_00_00000; // []
L[1072] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1073] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1074] = 9'b00_00_00000; // []
L[1075] = 9'b00_00_00000; // []
L[1076] = 9'b10_01_00110; // ALU()->[A0]
L[1077] = 9'b00_00_00000; // []
L[1078] = 9'b00_00_00000; // []
L[1079] = 9'b00_00_00000; // []
L[1080] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1081] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1082] = 9'b00_00_00000; // []
L[1083] = 9'b00_00_00000; // []
L[1084] = 9'b10_01_00110; // ALU()->[A0]
L[1085] = 9'b00_00_00000; // []
L[1086] = 9'b00_00_00000; // []
L[1087] = 9'b00_00_00000; // []
L[1088] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1089] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1090] = 9'b00_00_00000; // []
L[1091] = 9'b00_00_00000; // []
L[1092] = 9'b00_00_00000; // []
L[1093] = 9'b00_00_00000; // []
L[1094] = 9'b00_00_00000; // []
L[1095] = 9'b00_00_00000; // []
L[1096] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1097] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1098] = 9'b00_00_00000; // []
L[1099] = 9'b00_00_00000; // []
L[1100] = 9'b00_00_00000; // []
L[1101] = 9'b00_00_00000; // []
L[1102] = 9'b00_00_00000; // []
L[1103] = 9'b00_00_00000; // []
L[1104] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1105] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1106] = 9'b00_00_00000; // []
L[1107] = 9'b00_00_00000; // []
L[1108] = 9'b00_00_00000; // []
L[1109] = 9'b00_00_00000; // []
L[1110] = 9'b00_00_00000; // []
L[1111] = 9'b00_00_00000; // []
L[1112] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1113] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1114] = 9'b00_00_00000; // []
L[1115] = 9'b00_00_00000; // []
L[1116] = 9'b00_00_00000; // []
L[1117] = 9'b00_00_00000; // []
L[1118] = 9'b00_00_00000; // []
L[1119] = 9'b00_00_00000; // []
L[1120] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1121] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1122] = 9'b11_00_00001; // [PC++]->AH
L[1123] = 9'b00_00_00000; // []
L[1124] = 9'b10_01_00110; // ALU()->[A0]
L[1125] = 9'b00_00_00000; // []
L[1126] = 9'b00_00_00000; // []
L[1127] = 9'b00_00_00000; // []
L[1128] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1129] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1130] = 9'b11_00_00001; // [PC++]->AH
L[1131] = 9'b00_00_00000; // []
L[1132] = 9'b10_01_00110; // ALU()->[A0]
L[1133] = 9'b00_00_00000; // []
L[1134] = 9'b00_00_00000; // []
L[1135] = 9'b00_00_00000; // []
L[1136] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1137] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1138] = 9'b11_00_00001; // [PC++]->AH
L[1139] = 9'b00_00_00000; // []
L[1140] = 9'b10_01_00110; // ALU()->[A0]
L[1141] = 9'b00_00_00000; // []
L[1142] = 9'b00_00_00000; // []
L[1143] = 9'b00_00_00000; // []
L[1144] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1145] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1146] = 9'b11_00_00001; // [PC++]->AH
L[1147] = 9'b00_00_00000; // []
L[1148] = 9'b10_01_00110; // ALU()->[A0]
L[1149] = 9'b00_00_00000; // []
L[1150] = 9'b00_00_00000; // []
L[1151] = 9'b00_00_00000; // []
L[1152] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1153] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1154] = 9'b11_00_10001; // PC+T->PC
L[1155] = 9'b00_00_00000; // []
L[1156] = 9'b10_00_00011; // ['NO-OP', '']
L[1157] = 9'b00_00_00000; // []
L[1158] = 9'b00_00_00000; // []
L[1159] = 9'b00_00_00000; // []
L[1160] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1161] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1162] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1163] = 9'b00_01_01100; // [A0]->AH,T+Y->AL
L[1164] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1165] = 9'b10_01_00110; // ALU()->[A0]
L[1166] = 9'b00_00_00000; // []
L[1167] = 9'b00_00_00000; // []
L[1168] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1169] = 9'b10_00_00011; // ['NO-OP', '']
L[1170] = 9'b00_00_00000; // []
L[1171] = 9'b00_00_00000; // []
L[1172] = 9'b00_00_00000; // []
L[1173] = 9'b00_00_00000; // []
L[1174] = 9'b00_00_00000; // []
L[1175] = 9'b00_00_00000; // []
L[1176] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1177] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1178] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1179] = 9'b00_01_01100; // [A0]->AH,T+Y->AL
L[1180] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1181] = 9'b10_01_00110; // ALU()->[A0]
L[1182] = 9'b00_00_00000; // []
L[1183] = 9'b00_00_00000; // []
L[1184] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1185] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1186] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1187] = 9'b00_00_00000; // []
L[1188] = 9'b10_01_00110; // ALU()->[A0]
L[1189] = 9'b00_00_00000; // []
L[1190] = 9'b00_00_00000; // []
L[1191] = 9'b00_00_00000; // []
L[1192] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1193] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1194] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1195] = 9'b00_00_00000; // []
L[1196] = 9'b10_01_00110; // ALU()->[A0]
L[1197] = 9'b00_00_00000; // []
L[1198] = 9'b00_00_00000; // []
L[1199] = 9'b00_00_00000; // []
L[1200] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1201] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1202] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1203] = 9'b00_00_00000; // []
L[1204] = 9'b10_01_00110; // ALU()->[A0]
L[1205] = 9'b00_00_00000; // []
L[1206] = 9'b00_00_00000; // []
L[1207] = 9'b00_00_00000; // []
L[1208] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1209] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1210] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1211] = 9'b00_00_00000; // []
L[1212] = 9'b10_01_00110; // ALU()->[A0]
L[1213] = 9'b00_00_00000; // []
L[1214] = 9'b00_00_00000; // []
L[1215] = 9'b00_00_00000; // []
L[1216] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1217] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1218] = 9'b00_00_00000; // []
L[1219] = 9'b00_00_00000; // []
L[1220] = 9'b00_00_00000; // []
L[1221] = 9'b00_00_00000; // []
L[1222] = 9'b00_00_00000; // []
L[1223] = 9'b00_00_00000; // []
L[1224] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1225] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1226] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1227] = 9'b00_00_00000; // []
L[1228] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1229] = 9'b10_01_00110; // ALU()->[A0]
L[1230] = 9'b00_00_00000; // []
L[1231] = 9'b00_00_00000; // []
L[1232] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1233] = 9'b10_00_10010; // 0->S
L[1234] = 9'b00_00_00000; // []
L[1235] = 9'b00_00_00000; // []
L[1236] = 9'b00_00_00000; // []
L[1237] = 9'b00_00_00000; // []
L[1238] = 9'b00_00_00000; // []
L[1239] = 9'b00_00_00000; // []
L[1240] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1241] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1242] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1243] = 9'b00_00_00000; // []
L[1244] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1245] = 9'b10_01_00110; // ALU()->[A0]
L[1246] = 9'b00_00_00000; // []
L[1247] = 9'b00_00_00000; // []
L[1248] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1249] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1250] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1251] = 9'b00_00_00000; // []
L[1252] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1253] = 9'b10_01_00110; // ALU()->[A0]
L[1254] = 9'b00_00_00000; // []
L[1255] = 9'b00_00_00000; // []
L[1256] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1257] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1258] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1259] = 9'b00_00_00000; // []
L[1260] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1261] = 9'b10_01_00110; // ALU()->[A0]
L[1262] = 9'b00_00_00000; // []
L[1263] = 9'b00_00_00000; // []
L[1264] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1265] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1266] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1267] = 9'b00_00_00000; // []
L[1268] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1269] = 9'b10_01_00110; // ALU()->[A0]
L[1270] = 9'b00_00_00000; // []
L[1271] = 9'b00_00_00000; // []
L[1272] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1273] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1274] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1275] = 9'b00_00_00000; // []
L[1276] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1277] = 9'b10_01_00110; // ALU()->[A0]
L[1278] = 9'b00_00_00000; // []
L[1279] = 9'b00_00_00000; // []
L[1280] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1281] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[1282] = 9'b00_00_00000; // []
L[1283] = 9'b00_00_00000; // []
L[1284] = 9'b00_00_00000; // []
L[1285] = 9'b00_00_00000; // []
L[1286] = 9'b00_00_00000; // []
L[1287] = 9'b00_00_00000; // []
L[1288] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1289] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1290] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[1291] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1292] = 9'b00_01_01011; // [A0]->AH,T->AL
L[1293] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1294] = 9'b00_00_00000; // []
L[1295] = 9'b00_00_00000; // []
L[1296] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1297] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[1298] = 9'b00_00_00000; // []
L[1299] = 9'b00_00_00000; // []
L[1300] = 9'b00_00_00000; // []
L[1301] = 9'b00_00_00000; // []
L[1302] = 9'b00_00_00000; // []
L[1303] = 9'b00_00_00000; // []
L[1304] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1305] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1306] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[1307] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1308] = 9'b00_01_01011; // [A0]->AH,T->AL
L[1309] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1310] = 9'b00_00_00000; // []
L[1311] = 9'b00_00_00000; // []
L[1312] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1313] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1314] = 9'b00_00_00000; // []
L[1315] = 9'b00_00_00000; // []
L[1316] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1317] = 9'b00_00_00000; // []
L[1318] = 9'b00_00_00000; // []
L[1319] = 9'b00_00_00000; // []
L[1320] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1321] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1322] = 9'b00_00_00000; // []
L[1323] = 9'b00_00_00000; // []
L[1324] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1325] = 9'b00_00_00000; // []
L[1326] = 9'b00_00_00000; // []
L[1327] = 9'b00_00_00000; // []
L[1328] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1329] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1330] = 9'b00_00_00000; // []
L[1331] = 9'b00_00_00000; // []
L[1332] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1333] = 9'b00_00_00000; // []
L[1334] = 9'b00_00_00000; // []
L[1335] = 9'b00_00_00000; // []
L[1336] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1337] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1338] = 9'b00_00_00000; // []
L[1339] = 9'b00_00_00000; // []
L[1340] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1341] = 9'b00_00_00000; // []
L[1342] = 9'b00_00_00000; // []
L[1343] = 9'b00_00_00000; // []
L[1344] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1345] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1346] = 9'b00_00_00000; // []
L[1347] = 9'b00_00_00000; // []
L[1348] = 9'b00_00_00000; // []
L[1349] = 9'b00_00_00000; // []
L[1350] = 9'b00_00_00000; // []
L[1351] = 9'b00_00_00000; // []
L[1352] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1353] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[1354] = 9'b00_00_00000; // []
L[1355] = 9'b00_00_00000; // []
L[1356] = 9'b00_00_00000; // []
L[1357] = 9'b00_00_00000; // []
L[1358] = 9'b00_00_00000; // []
L[1359] = 9'b00_00_00000; // []
L[1360] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1361] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1362] = 9'b00_00_00000; // []
L[1363] = 9'b00_00_00000; // []
L[1364] = 9'b00_00_00000; // []
L[1365] = 9'b00_00_00000; // []
L[1366] = 9'b00_00_00000; // []
L[1367] = 9'b00_00_00000; // []
L[1368] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1369] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1370] = 9'b00_00_00000; // []
L[1371] = 9'b00_00_00000; // []
L[1372] = 9'b00_00_00000; // []
L[1373] = 9'b00_00_00000; // []
L[1374] = 9'b00_00_00000; // []
L[1375] = 9'b00_00_00000; // []
L[1376] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1377] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1378] = 9'b11_00_00001; // [PC++]->AH
L[1379] = 9'b00_00_00000; // []
L[1380] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1381] = 9'b00_00_00000; // []
L[1382] = 9'b00_00_00000; // []
L[1383] = 9'b00_00_00000; // []
L[1384] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1385] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1386] = 9'b11_00_00001; // [PC++]->AH
L[1387] = 9'b00_00_00000; // []
L[1388] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1389] = 9'b00_00_00000; // []
L[1390] = 9'b00_00_00000; // []
L[1391] = 9'b00_00_00000; // []
L[1392] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1393] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1394] = 9'b11_00_00001; // [PC++]->AH
L[1395] = 9'b00_00_00000; // []
L[1396] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1397] = 9'b00_00_00000; // []
L[1398] = 9'b00_00_00000; // []
L[1399] = 9'b00_00_00000; // []
L[1400] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1401] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1402] = 9'b11_00_00001; // [PC++]->AH
L[1403] = 9'b00_00_00000; // []
L[1404] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1405] = 9'b00_00_00000; // []
L[1406] = 9'b00_00_00000; // []
L[1407] = 9'b00_00_00000; // []
L[1408] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1409] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1410] = 9'b11_00_10001; // PC+T->PC
L[1411] = 9'b00_00_00000; // []
L[1412] = 9'b10_00_00011; // ['NO-OP', '']
L[1413] = 9'b00_00_00000; // []
L[1414] = 9'b00_00_00000; // []
L[1415] = 9'b00_00_00000; // []
L[1416] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1417] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1418] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1419] = 9'b01_01_01100; // [A0]->AH,T+Y->AL
L[1420] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1421] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1422] = 9'b00_00_00000; // []
L[1423] = 9'b00_00_00000; // []
L[1424] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1425] = 9'b10_00_00011; // ['NO-OP', '']
L[1426] = 9'b00_00_00000; // []
L[1427] = 9'b00_00_00000; // []
L[1428] = 9'b00_00_00000; // []
L[1429] = 9'b00_00_00000; // []
L[1430] = 9'b00_00_00000; // []
L[1431] = 9'b00_00_00000; // []
L[1432] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1433] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1434] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1435] = 9'b01_01_01100; // [A0]->AH,T+Y->AL
L[1436] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1437] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1438] = 9'b00_00_00000; // []
L[1439] = 9'b00_00_00000; // []
L[1440] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1441] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1442] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1443] = 9'b00_00_00000; // []
L[1444] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1445] = 9'b00_00_00000; // []
L[1446] = 9'b00_00_00000; // []
L[1447] = 9'b00_00_00000; // []
L[1448] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1449] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1450] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1451] = 9'b00_00_00000; // []
L[1452] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1453] = 9'b00_00_00000; // []
L[1454] = 9'b00_00_00000; // []
L[1455] = 9'b00_00_00000; // []
L[1456] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1457] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1458] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1459] = 9'b00_00_00000; // []
L[1460] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1461] = 9'b00_00_00000; // []
L[1462] = 9'b00_00_00000; // []
L[1463] = 9'b00_00_00000; // []
L[1464] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1465] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1466] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1467] = 9'b00_00_00000; // []
L[1468] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1469] = 9'b00_00_00000; // []
L[1470] = 9'b00_00_00000; // []
L[1471] = 9'b00_00_00000; // []
L[1472] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1473] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1474] = 9'b00_00_00000; // []
L[1475] = 9'b00_00_00000; // []
L[1476] = 9'b00_00_00000; // []
L[1477] = 9'b00_00_00000; // []
L[1478] = 9'b00_00_00000; // []
L[1479] = 9'b00_00_00000; // []
L[1480] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1481] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1482] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1483] = 9'b00_00_00000; // []
L[1484] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1485] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1486] = 9'b00_00_00000; // []
L[1487] = 9'b00_00_00000; // []
L[1488] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1489] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1490] = 9'b00_00_00000; // []
L[1491] = 9'b00_00_00000; // []
L[1492] = 9'b00_00_00000; // []
L[1493] = 9'b00_00_00000; // []
L[1494] = 9'b00_00_00000; // []
L[1495] = 9'b00_00_00000; // []
L[1496] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1497] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1498] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1499] = 9'b00_00_00000; // []
L[1500] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1501] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1502] = 9'b00_00_00000; // []
L[1503] = 9'b00_00_00000; // []
L[1504] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1505] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1506] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1507] = 9'b00_00_00000; // []
L[1508] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1509] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1510] = 9'b00_00_00000; // []
L[1511] = 9'b00_00_00000; // []
L[1512] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1513] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1514] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1515] = 9'b00_00_00000; // []
L[1516] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1517] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1518] = 9'b00_00_00000; // []
L[1519] = 9'b00_00_00000; // []
L[1520] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1521] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1522] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1523] = 9'b00_00_00000; // []
L[1524] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1525] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1526] = 9'b00_00_00000; // []
L[1527] = 9'b00_00_00000; // []
L[1528] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1529] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1530] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1531] = 9'b00_00_00000; // []
L[1532] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1533] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1534] = 9'b00_00_00000; // []
L[1535] = 9'b00_00_00000; // []
L[1536] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1537] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[1538] = 9'b00_00_00000; // []
L[1539] = 9'b00_00_00000; // []
L[1540] = 9'b00_00_00000; // []
L[1541] = 9'b00_00_00000; // []
L[1542] = 9'b00_00_00000; // []
L[1543] = 9'b00_00_00000; // []
L[1544] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1545] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1546] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[1547] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1548] = 9'b00_01_01011; // [A0]->AH,T->AL
L[1549] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1550] = 9'b00_00_00000; // []
L[1551] = 9'b00_00_00000; // []
L[1552] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1553] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1554] = 9'b00_00_00000; // []
L[1555] = 9'b00_00_00000; // []
L[1556] = 9'b00_00_00000; // []
L[1557] = 9'b00_00_00000; // []
L[1558] = 9'b00_00_00000; // []
L[1559] = 9'b00_00_00000; // []
L[1560] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1561] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1562] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[1563] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1564] = 9'b00_01_01011; // [A0]->AH,T->AL
L[1565] = 9'b00_01_00011; // [A0]->T
L[1566] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1567] = 9'b10_01_00101; // T->[A0]
L[1568] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1569] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1570] = 9'b00_00_00000; // []
L[1571] = 9'b00_00_00000; // []
L[1572] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1573] = 9'b00_00_00000; // []
L[1574] = 9'b00_00_00000; // []
L[1575] = 9'b00_00_00000; // []
L[1576] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1577] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1578] = 9'b00_00_00000; // []
L[1579] = 9'b00_00_00000; // []
L[1580] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1581] = 9'b00_00_00000; // []
L[1582] = 9'b00_00_00000; // []
L[1583] = 9'b00_00_00000; // []
L[1584] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1585] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1586] = 9'b00_00_00000; // []
L[1587] = 9'b00_00_00000; // []
L[1588] = 9'b00_01_00011; // [A0]->T
L[1589] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1590] = 9'b10_01_00101; // T->[A0]
L[1591] = 9'b00_00_00000; // []
L[1592] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1593] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1594] = 9'b00_00_00000; // []
L[1595] = 9'b00_00_00000; // []
L[1596] = 9'b00_01_00011; // [A0]->T
L[1597] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1598] = 9'b10_01_00101; // T->[A0]
L[1599] = 9'b00_00_00000; // []
L[1600] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1601] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1602] = 9'b00_00_00000; // []
L[1603] = 9'b00_00_00000; // []
L[1604] = 9'b00_00_00000; // []
L[1605] = 9'b00_00_00000; // []
L[1606] = 9'b00_00_00000; // []
L[1607] = 9'b00_00_00000; // []
L[1608] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1609] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[1610] = 9'b00_00_00000; // []
L[1611] = 9'b00_00_00000; // []
L[1612] = 9'b00_00_00000; // []
L[1613] = 9'b00_00_00000; // []
L[1614] = 9'b00_00_00000; // []
L[1615] = 9'b00_00_00000; // []
L[1616] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1617] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1618] = 9'b00_00_00000; // []
L[1619] = 9'b00_00_00000; // []
L[1620] = 9'b00_00_00000; // []
L[1621] = 9'b00_00_00000; // []
L[1622] = 9'b00_00_00000; // []
L[1623] = 9'b00_00_00000; // []
L[1624] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1625] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1626] = 9'b00_00_00000; // []
L[1627] = 9'b00_00_00000; // []
L[1628] = 9'b00_00_00000; // []
L[1629] = 9'b00_00_00000; // []
L[1630] = 9'b00_00_00000; // []
L[1631] = 9'b00_00_00000; // []
L[1632] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1633] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1634] = 9'b11_00_00001; // [PC++]->AH
L[1635] = 9'b00_00_00000; // []
L[1636] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1637] = 9'b00_00_00000; // []
L[1638] = 9'b00_00_00000; // []
L[1639] = 9'b00_00_00000; // []
L[1640] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1641] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1642] = 9'b11_00_00001; // [PC++]->AH
L[1643] = 9'b00_00_00000; // []
L[1644] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1645] = 9'b00_00_00000; // []
L[1646] = 9'b00_00_00000; // []
L[1647] = 9'b00_00_00000; // []
L[1648] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1649] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1650] = 9'b11_00_00001; // [PC++]->AH
L[1651] = 9'b00_00_00000; // []
L[1652] = 9'b00_01_00011; // [A0]->T
L[1653] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1654] = 9'b10_01_00101; // T->[A0]
L[1655] = 9'b00_00_00000; // []
L[1656] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1657] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1658] = 9'b11_00_00001; // [PC++]->AH
L[1659] = 9'b00_00_00000; // []
L[1660] = 9'b00_01_00011; // [A0]->T
L[1661] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1662] = 9'b10_01_00101; // T->[A0]
L[1663] = 9'b00_00_00000; // []
L[1664] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1665] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1666] = 9'b11_00_10001; // PC+T->PC
L[1667] = 9'b00_00_00000; // []
L[1668] = 9'b10_00_00011; // ['NO-OP', '']
L[1669] = 9'b00_00_00000; // []
L[1670] = 9'b00_00_00000; // []
L[1671] = 9'b00_00_00000; // []
L[1672] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1673] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1674] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1675] = 9'b01_01_01100; // [A0]->AH,T+Y->AL
L[1676] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1677] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1678] = 9'b00_00_00000; // []
L[1679] = 9'b00_00_00000; // []
L[1680] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1681] = 9'b10_00_00011; // ['NO-OP', '']
L[1682] = 9'b00_00_00000; // []
L[1683] = 9'b00_00_00000; // []
L[1684] = 9'b00_00_00000; // []
L[1685] = 9'b00_00_00000; // []
L[1686] = 9'b00_00_00000; // []
L[1687] = 9'b00_00_00000; // []
L[1688] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1689] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1690] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1691] = 9'b00_01_01100; // [A0]->AH,T+Y->AL
L[1692] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1693] = 9'b00_01_00011; // [A0]->T
L[1694] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1695] = 9'b10_01_00101; // T->[A0]
L[1696] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1697] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1698] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1699] = 9'b00_00_00000; // []
L[1700] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[1701] = 9'b00_00_00000; // []
L[1702] = 9'b00_00_00000; // []
L[1703] = 9'b00_00_00000; // []
L[1704] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1705] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1706] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1707] = 9'b00_00_00000; // []
L[1708] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1709] = 9'b00_00_00000; // []
L[1710] = 9'b00_00_00000; // []
L[1711] = 9'b00_00_00000; // []
L[1712] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1713] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1714] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1715] = 9'b00_00_00000; // []
L[1716] = 9'b00_01_00011; // [A0]->T
L[1717] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1718] = 9'b10_01_00101; // T->[A0]
L[1719] = 9'b00_00_00000; // []
L[1720] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1721] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1722] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1723] = 9'b00_00_00000; // []
L[1724] = 9'b00_01_00011; // [A0]->T
L[1725] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1726] = 9'b10_01_00101; // T->[A0]
L[1727] = 9'b00_00_00000; // []
L[1728] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1729] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1730] = 9'b00_00_00000; // []
L[1731] = 9'b00_00_00000; // []
L[1732] = 9'b00_00_00000; // []
L[1733] = 9'b00_00_00000; // []
L[1734] = 9'b00_00_00000; // []
L[1735] = 9'b00_00_00000; // []
L[1736] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1737] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1738] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1739] = 9'b00_00_00000; // []
L[1740] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1741] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1742] = 9'b00_00_00000; // []
L[1743] = 9'b00_00_00000; // []
L[1744] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1745] = 9'b10_00_00011; // ['NO-OP', '']
L[1746] = 9'b00_00_00000; // []
L[1747] = 9'b00_00_00000; // []
L[1748] = 9'b00_00_00000; // []
L[1749] = 9'b00_00_00000; // []
L[1750] = 9'b00_00_00000; // []
L[1751] = 9'b00_00_00000; // []
L[1752] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1753] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1754] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1755] = 9'b00_00_00000; // []
L[1756] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1757] = 9'b00_01_00011; // [A0]->T
L[1758] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1759] = 9'b10_01_00101; // T->[A0]
L[1760] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1761] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1762] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1763] = 9'b00_00_00000; // []
L[1764] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1765] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[1766] = 9'b00_00_00000; // []
L[1767] = 9'b00_00_00000; // []
L[1768] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1769] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1770] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1771] = 9'b00_00_00000; // []
L[1772] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1773] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1774] = 9'b00_00_00000; // []
L[1775] = 9'b00_00_00000; // []
L[1776] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1777] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1778] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1779] = 9'b00_00_00000; // []
L[1780] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1781] = 9'b00_01_00011; // [A0]->T
L[1782] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1783] = 9'b10_01_00101; // T->[A0]
L[1784] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1785] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1786] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1787] = 9'b00_00_00000; // []
L[1788] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1789] = 9'b00_01_00011; // [A0]->T
L[1790] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1791] = 9'b10_01_00101; // T->[A0]
L[1792] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1793] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[1794] = 9'b00_00_00000; // []
L[1795] = 9'b00_00_00000; // []
L[1796] = 9'b00_00_00000; // []
L[1797] = 9'b00_00_00000; // []
L[1798] = 9'b00_00_00000; // []
L[1799] = 9'b00_00_00000; // []
L[1800] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1801] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1802] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[1803] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1804] = 9'b00_01_01011; // [A0]->AH,T->AL
L[1805] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1806] = 9'b00_00_00000; // []
L[1807] = 9'b00_00_00000; // []
L[1808] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1809] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1810] = 9'b00_00_00000; // []
L[1811] = 9'b00_00_00000; // []
L[1812] = 9'b00_00_00000; // []
L[1813] = 9'b00_00_00000; // []
L[1814] = 9'b00_00_00000; // []
L[1815] = 9'b00_00_00000; // []
L[1816] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1817] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1818] = 9'b00_01_00111; // [A0]->?,AL+0->AL
L[1819] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1820] = 9'b00_01_01011; // [A0]->AH,T->AL
L[1821] = 9'b00_01_00011; // [A0]->T
L[1822] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1823] = 9'b10_01_00101; // T->[A0]
L[1824] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1825] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1826] = 9'b00_00_00000; // []
L[1827] = 9'b00_00_00000; // []
L[1828] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1829] = 9'b00_00_00000; // []
L[1830] = 9'b00_00_00000; // []
L[1831] = 9'b00_00_00000; // []
L[1832] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1833] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1834] = 9'b00_00_00000; // []
L[1835] = 9'b00_00_00000; // []
L[1836] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1837] = 9'b00_00_00000; // []
L[1838] = 9'b00_00_00000; // []
L[1839] = 9'b00_00_00000; // []
L[1840] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1841] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1842] = 9'b00_00_00000; // []
L[1843] = 9'b00_00_00000; // []
L[1844] = 9'b00_01_00011; // [A0]->T
L[1845] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1846] = 9'b10_01_00101; // T->[A0]
L[1847] = 9'b00_00_00000; // []
L[1848] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1849] = 9'b11_00_00000; // ['[PC++]->AL', '[PC++]->T']
L[1850] = 9'b00_00_00000; // []
L[1851] = 9'b00_00_00000; // []
L[1852] = 9'b00_01_00011; // [A0]->T
L[1853] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1854] = 9'b10_01_00101; // T->[A0]
L[1855] = 9'b00_00_00000; // []
L[1856] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1857] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1858] = 9'b00_00_00000; // []
L[1859] = 9'b00_00_00000; // []
L[1860] = 9'b00_00_00000; // []
L[1861] = 9'b00_00_00000; // []
L[1862] = 9'b00_00_00000; // []
L[1863] = 9'b00_00_00000; // []
L[1864] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1865] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[1866] = 9'b00_00_00000; // []
L[1867] = 9'b00_00_00000; // []
L[1868] = 9'b00_00_00000; // []
L[1869] = 9'b00_00_00000; // []
L[1870] = 9'b00_00_00000; // []
L[1871] = 9'b00_00_00000; // []
L[1872] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1873] = 9'b10_00_00011; // ['NO-OP', '']
L[1874] = 9'b00_00_00000; // []
L[1875] = 9'b00_00_00000; // []
L[1876] = 9'b00_00_00000; // []
L[1877] = 9'b00_00_00000; // []
L[1878] = 9'b00_00_00000; // []
L[1879] = 9'b00_00_00000; // []
L[1880] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1881] = 9'b10_00_01101; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
L[1882] = 9'b00_00_00000; // []
L[1883] = 9'b00_00_00000; // []
L[1884] = 9'b00_00_00000; // []
L[1885] = 9'b00_00_00000; // []
L[1886] = 9'b00_00_00000; // []
L[1887] = 9'b00_00_00000; // []
L[1888] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1889] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1890] = 9'b11_00_00001; // [PC++]->AH
L[1891] = 9'b00_00_00000; // []
L[1892] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1893] = 9'b00_00_00000; // []
L[1894] = 9'b00_00_00000; // []
L[1895] = 9'b00_00_00000; // []
L[1896] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1897] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1898] = 9'b11_00_00001; // [PC++]->AH
L[1899] = 9'b00_00_00000; // []
L[1900] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1901] = 9'b00_00_00000; // []
L[1902] = 9'b00_00_00000; // []
L[1903] = 9'b00_00_00000; // []
L[1904] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1905] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1906] = 9'b11_00_00001; // [PC++]->AH
L[1907] = 9'b00_00_00000; // []
L[1908] = 9'b00_01_00011; // [A0]->T
L[1909] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1910] = 9'b10_01_00101; // T->[A0]
L[1911] = 9'b00_00_00000; // []
L[1912] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1913] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1914] = 9'b11_00_00001; // [PC++]->AH
L[1915] = 9'b00_00_00000; // []
L[1916] = 9'b00_01_00011; // [A0]->T
L[1917] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1918] = 9'b10_01_00101; // T->[A0]
L[1919] = 9'b00_00_00000; // []
L[1920] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1921] = 9'b10_00_00000; // ['[PC++]->?', 'PC+1->PC', '']
L[1922] = 9'b11_00_10001; // PC+T->PC
L[1923] = 9'b00_00_00000; // []
L[1924] = 9'b10_00_00011; // ['NO-OP', '']
L[1925] = 9'b00_00_00000; // []
L[1926] = 9'b00_00_00000; // []
L[1927] = 9'b00_00_00000; // []
L[1928] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1929] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1930] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1931] = 9'b01_01_01100; // [A0]->AH,T+Y->AL
L[1932] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1933] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1934] = 9'b00_00_00000; // []
L[1935] = 9'b00_00_00000; // []
L[1936] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1937] = 9'b10_00_00011; // ['NO-OP', '']
L[1938] = 9'b00_00_00000; // []
L[1939] = 9'b00_00_00000; // []
L[1940] = 9'b00_00_00000; // []
L[1941] = 9'b00_00_00000; // []
L[1942] = 9'b00_00_00000; // []
L[1943] = 9'b00_00_00000; // []
L[1944] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1945] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1946] = 9'b00_01_01010; // [A0]->T,AL+1->AL
L[1947] = 9'b00_01_01100; // [A0]->AH,T+Y->AL
L[1948] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1949] = 9'b00_01_00011; // [A0]->T
L[1950] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1951] = 9'b10_01_00101; // T->[A0]
L[1952] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1953] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1954] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1955] = 9'b00_00_00000; // []
L[1956] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[1957] = 9'b00_00_00000; // []
L[1958] = 9'b00_00_00000; // []
L[1959] = 9'b00_00_00000; // []
L[1960] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1961] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1962] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1963] = 9'b00_00_00000; // []
L[1964] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1965] = 9'b00_00_00000; // []
L[1966] = 9'b00_00_00000; // []
L[1967] = 9'b00_00_00000; // []
L[1968] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1969] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1970] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1971] = 9'b00_00_00000; // []
L[1972] = 9'b00_01_00011; // [A0]->T
L[1973] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1974] = 9'b10_01_00101; // T->[A0]
L[1975] = 9'b00_00_00000; // []
L[1976] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1977] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1978] = 9'b11_01_00111; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL']
L[1979] = 9'b00_00_00000; // []
L[1980] = 9'b00_01_00011; // [A0]->T
L[1981] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[1982] = 9'b10_01_00101; // T->[A0]
L[1983] = 9'b00_00_00000; // []
L[1984] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1985] = 9'b10_00_00010; // ['[PC]->,ALU()->A', 'Setappropriateflags', 'ALU()->0,Y', 'ALU()->A']
L[1986] = 9'b00_00_00000; // []
L[1987] = 9'b00_00_00000; // []
L[1988] = 9'b00_00_00000; // []
L[1989] = 9'b00_00_00000; // []
L[1990] = 9'b00_00_00000; // []
L[1991] = 9'b00_00_00000; // []
L[1992] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1993] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[1994] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[1995] = 9'b00_00_00000; // []
L[1996] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[1997] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[1998] = 9'b00_00_00000; // []
L[1999] = 9'b00_00_00000; // []
L[2000] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2001] = 9'b10_00_00011; // ['NO-OP', '']
L[2002] = 9'b00_00_00000; // []
L[2003] = 9'b00_00_00000; // []
L[2004] = 9'b00_00_00000; // []
L[2005] = 9'b00_00_00000; // []
L[2006] = 9'b00_00_00000; // []
L[2007] = 9'b00_00_00000; // []
L[2008] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2009] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2010] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[2011] = 9'b00_00_00000; // []
L[2012] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[2013] = 9'b00_01_00011; // [A0]->T
L[2014] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[2015] = 9'b10_01_00101; // T->[A0]
L[2016] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2017] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2018] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[2019] = 9'b00_00_00000; // []
L[2020] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[2021] = 9'b10_01_00011; // ['ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->']
L[2022] = 9'b00_00_00000; // []
L[2023] = 9'b00_00_00000; // []
L[2024] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2025] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2026] = 9'b01_00_01000; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[2027] = 9'b00_00_00000; // []
L[2028] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[2029] = 9'b10_01_00010; // ['ALU([A0])->A', 'ALU([A0])->?']
L[2030] = 9'b00_00_00000; // []
L[2031] = 9'b00_00_00000; // []
L[2032] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2033] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2034] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[2035] = 9'b00_00_00000; // []
L[2036] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[2037] = 9'b00_01_00011; // [A0]->T
L[2038] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[2039] = 9'b10_01_00101; // T->[A0]
L[2040] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2041] = 9'b00_00_00000; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T']
L[2042] = 9'b11_00_01000; // ['[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+Y->AL']
L[2043] = 9'b00_00_00000; // []
L[2044] = 9'b00_01_01001; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
L[2045] = 9'b00_01_00011; // [A0]->T
L[2046] = 9'b00_01_00100; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
L[2047] = 9'b10_01_00101; // T->[A0]
  end  
  always @(posedge clk) if (reset) begin
    M <= 0; // Stupid XILINX inferral only allows 0 as reset value.
  end else if (ce) begin
    M <= L[{IR, State}];    
  end
endmodule

module MicroCodeTable(input clk, input ce, input reset, input [7:0] IR, input [2:0] State, output [37:0] Mout);
  wire [8:0] M;
  MicroCodeTableInner inner(clk, ce, reset, IR, State, M);
  reg [14:0] A[0:31];
  reg [18:0] B[0:255];
  initial begin
A[0] = 15'b_10__0_10101_000_01_00; // ['[PC++]', '[PC++]->AL', '[PC++]->?', '[PC++]->T', 'PC+1->PC', '']
A[1] = 15'b_00__0_00011_000_01_00; // [PC++]->AH
A[2] = 15'b_00__1_00000_000_00_00; // ['ALU([A0])->A', 'ALU([A0])->?', '[PC]->,ALU()->A', 'Setappropriateflags', 'ALU([SP])->A', '[SP]->P', 'ALU()->0,Y', 'ALU()->A']
A[3] = 15'b_10__0_00000_000_00_00; // ['[A0]->T', 'ALU([A0])->?', 'ALU([A0])->A', 'ALU([A0])->', '[PC]->', 'NO-OP', '[VECT]->T', '']
A[4] = 15'b_11__1_00000_100_00_00; // ['T->[A0],ALU(T)->T', 'T->[A0],ALU(T)->T:A']
A[5] = 15'b_00__0_00000_100_00_00; // T->[A0]
A[6] = 15'b_00__0_00000_101_00_00; // ALU()->[A0]
A[7] = 15'b_00__0_10000_000_00_00; // ['[A0]->?,AL+0->AL', '[A0]->?,AL+0/Y->AL', 'KEEP_AC']
A[8] = 15'b_00__0_10011_000_01_00; // ['[PC++]->AH,AL+0/Y->AL', '[PC++]->AH,AL+0->AL', '[PC++]->AH,AL+Y->AL']
A[9] = 15'b_10__0_00010_000_00_00; // ['[A0]->?,AH+FI0->AH', '[A0]->T,AH+FI0->AH']
A[10] = 15'b_10__0_11000_000_00_00; // [A0]->T,AL+1->AL
A[11] = 15'b_00__0_11111_000_00_00; // [A0]->AH,T->AL
A[12] = 15'b_00__0_10011_000_00_00; // [A0]->AH,T+Y->AL
A[13] = 15'b_00__1_00000_000_01_00; // ['ALU([PC++])->A', 'ALU([PC++])->?', 'ALU([PC++])->Reg']
A[14] = 15'b_00__0_00000_101_00_11; // ALU(A)->[SP--]
A[15] = 15'b_00__0_00000_110_00_11; // P->[SP--]
A[16] = 15'b_10__0_00000_000_00_10; // ['SP++', 'SP+1->SP', '[SP]->T,SP+1->SP']
A[17] = 15'b_00__0_00000_000_11_00; // PC+T->PC
A[18] = 15'b_00__0_00000_000_00_01; // 0->S
A[19] = 15'b_00__0_00000_000_10_00; // ['[PC]:T->PC', '[A0]:T->PC', '[VECT]:T->PC', '[SP]:T->PC']
A[20] = 15'b_00__0_00000_111_00_11; // ['PCH->[SP--]', 'PCL->[SP--],', 'PCH->[SP--](KEEPAC)', 'PCL->[SP--](KEEPAC)']
A[21] = 15'b_00__1_00000_110_00_11; // P->[SP--]
A[22] = 15'b_00__1_00000_000_00_10; // [SP]->P,SP+1->SP
A[23] = 15'b_00__0_00000_000_00_00; // []
A[24] = 15'b_00__0_00000_000_00_00; // []
A[25] = 15'b_00__0_00000_000_00_00; // []
A[26] = 15'b_00__0_00000_000_00_00; // []
A[27] = 15'b_00__0_00000_000_00_00; // []
A[28] = 15'b_00__0_00000_000_00_00; // []
A[29] = 15'b_00__0_00000_000_00_00; // []
A[30] = 15'b_00__0_00000_000_00_00; // []
A[31] = 15'b_00__0_00000_000_00_00; // []
B[0] = 19'b00000000000_000_00_010;
B[32] = 19'b00000000000_000_00_000;
B[64] = 19'b00000000000_000_00_100;
B[96] = 19'b00000000000_000_00_000;
B[128] = 19'b01101001000_000_00_000;
B[160] = 19'b00001001000_100_00_001;
B[192] = 19'b01001001100_000_00_001;
B[224] = 19'b10001001100_000_00_001;
B[1] = 19'b00001000001_010_00_001;
B[33] = 19'b00001000011_010_00_001;
B[65] = 19'b00001000101_010_00_001;
B[97] = 19'b00001000111_010_00_001;
B[129] = 19'b00101001001_000_00_000;
B[161] = 19'b00001001001_010_00_001;
B[193] = 19'b00001001101_000_00_001;
B[225] = 19'b00001001111_010_00_001;
B[2] = 19'b00010001000_000_00_001;
B[34] = 19'b00010011000_000_00_001;
B[66] = 19'b00010101000_000_00_001;
B[98] = 19'b00010111000_000_00_001;
B[130] = 19'b10101001000_000_00_000;
B[162] = 19'b00001001000_001_00_001;
B[194] = 19'b00011101000_000_00_001;
B[226] = 19'b00011111000_000_00_001;
B[3] = 19'b00010000001_010_00_001;
B[35] = 19'b00010010011_010_00_001;
B[67] = 19'b00010100101_010_00_001;
B[99] = 19'b00010110111_010_00_001;
B[131] = 19'b11101001001_000_00_000;
B[163] = 19'b00001001001_011_00_001;
B[195] = 19'b00011101101_000_00_001;
B[227] = 19'b00011111111_010_00_001;
B[4] = 19'b00001000000_000_00_000;
B[36] = 19'b00001000010_000_00_001;
B[68] = 19'b00001000100_000_00_000;
B[100] = 19'b00001000110_000_00_000;
B[132] = 19'b01101001000_000_00_000;
B[164] = 19'b00001001000_100_00_001;
B[196] = 19'b01001001100_000_00_001;
B[228] = 19'b10001001100_000_00_001;
B[5] = 19'b00001000001_010_00_001;
B[37] = 19'b00001000011_010_00_001;
B[69] = 19'b00001000101_010_00_001;
B[101] = 19'b00001000111_010_00_001;
B[133] = 19'b00101001001_000_00_000;
B[165] = 19'b00001001001_010_00_001;
B[197] = 19'b00001001101_000_00_001;
B[229] = 19'b00001001111_010_00_001;
B[6] = 19'b00010001000_000_00_001;
B[38] = 19'b00010011000_000_00_001;
B[70] = 19'b00010101000_000_00_001;
B[102] = 19'b00010111000_000_00_001;
B[134] = 19'b10101001000_000_00_000;
B[166] = 19'b00001001000_001_00_001;
B[198] = 19'b00011101000_000_00_001;
B[230] = 19'b00011111000_000_00_001;
B[7] = 19'b00010000001_010_00_001;
B[39] = 19'b00010010011_010_00_001;
B[71] = 19'b00010100101_010_00_001;
B[103] = 19'b00010110111_010_00_001;
B[135] = 19'b11101001001_000_00_000;
B[167] = 19'b00001001001_011_00_001;
B[199] = 19'b00011101101_000_00_001;
B[231] = 19'b00011111111_010_00_001;
B[8] = 19'b00000000000_000_00_000;
B[40] = 19'b00000000000_000_00_100;
B[72] = 19'b00101001000_000_00_000;
B[104] = 19'b00001001000_010_00_001;
B[136] = 19'b01101101000_100_00_001;
B[168] = 19'b00101001000_100_00_001;
B[200] = 19'b01101111000_100_00_001;
B[232] = 19'b10101111000_001_00_001;
B[9] = 19'b00001000001_010_00_001;
B[41] = 19'b00001000011_010_00_001;
B[73] = 19'b00001000101_010_00_001;
B[105] = 19'b00001000111_010_00_001;
B[137] = 19'b00101001001_000_00_000;
B[169] = 19'b00001001001_010_00_001;
B[201] = 19'b00001001101_000_00_001;
B[233] = 19'b00001001111_010_00_001;
B[10] = 19'b00100001000_010_00_001;
B[42] = 19'b00100011000_010_00_001;
B[74] = 19'b00100101000_010_00_001;
B[106] = 19'b00100111000_010_00_001;
B[138] = 19'b10101001000_010_00_001;
B[170] = 19'b00101001000_001_00_001;
B[202] = 19'b10101101000_001_00_001;
B[234] = 19'b00011111000_000_00_001;
B[11] = 19'b00001000001_010_00_001;
B[43] = 19'b00001000011_010_00_001;
B[75] = 19'b00001000101_010_00_001;
B[107] = 19'b00001000111_010_00_001;
B[139] = 19'b11101001001_000_00_000;
B[171] = 19'b00001001001_011_00_001;
B[203] = 19'b00001001101_000_00_001;
B[235] = 19'b00001001111_010_00_001;
B[12] = 19'b00001000000_000_00_000;
B[44] = 19'b00001000010_000_00_001;
B[76] = 19'b00000000000_000_00_001;
B[108] = 19'b00000000000_000_00_001;
B[140] = 19'b01101001000_000_00_000;
B[172] = 19'b00001001000_100_00_001;
B[204] = 19'b01001001100_000_00_001;
B[236] = 19'b10001001100_000_00_001;
B[13] = 19'b00001000001_010_00_001;
B[45] = 19'b00001000011_010_00_001;
B[77] = 19'b00001000101_010_00_001;
B[109] = 19'b00001000111_010_00_001;
B[141] = 19'b00101001001_000_00_000;
B[173] = 19'b00001001001_010_00_001;
B[205] = 19'b00001001101_000_00_001;
B[237] = 19'b00001001111_010_00_001;
B[14] = 19'b00010001000_000_00_001;
B[46] = 19'b00010011000_000_00_001;
B[78] = 19'b00010101000_000_00_001;
B[110] = 19'b00010111000_000_00_001;
B[142] = 19'b10101001000_000_00_000;
B[174] = 19'b00001001000_001_00_001;
B[206] = 19'b00011101000_000_00_001;
B[238] = 19'b00011111000_000_00_001;
B[15] = 19'b00010000001_010_00_001;
B[47] = 19'b00010010011_010_00_001;
B[79] = 19'b00010100101_010_00_001;
B[111] = 19'b00010110111_010_00_001;
B[143] = 19'b11101001001_000_00_000;
B[175] = 19'b00001001001_011_00_001;
B[207] = 19'b00011101101_000_00_001;
B[239] = 19'b00011111111_010_00_001;
B[16] = 19'b00000000000_000_11_000;
B[48] = 19'b00000000000_000_11_000;
B[80] = 19'b00000000000_000_11_000;
B[112] = 19'b00000000000_000_11_000;
B[144] = 19'b01101001000_000_11_000;
B[176] = 19'b00001001000_000_11_000;
B[208] = 19'b00000000000_000_11_000;
B[240] = 19'b00000000000_000_11_000;
B[17] = 19'b00001000001_010_11_001;
B[49] = 19'b00001000011_010_11_001;
B[81] = 19'b00001000101_010_11_001;
B[113] = 19'b00001000111_010_11_001;
B[145] = 19'b00101001001_000_11_000;
B[177] = 19'b00001001001_010_11_001;
B[209] = 19'b00001001101_000_11_001;
B[241] = 19'b00001001111_010_11_001;
B[18] = 19'b00010001000_000_11_001;
B[50] = 19'b00010011000_000_11_001;
B[82] = 19'b00010101000_000_11_001;
B[114] = 19'b00010111000_000_11_001;
B[146] = 19'b10101001000_000_11_000;
B[178] = 19'b00001001000_000_11_000;
B[210] = 19'b00011101000_000_11_001;
B[242] = 19'b00011111000_000_11_001;
B[19] = 19'b00010000001_010_11_001;
B[51] = 19'b00010010011_010_11_001;
B[83] = 19'b00010100101_010_11_001;
B[115] = 19'b00010110111_010_11_001;
B[147] = 19'b11101001001_000_11_000;
B[179] = 19'b00001001001_011_11_001;
B[211] = 19'b00011101101_000_11_001;
B[243] = 19'b00011111111_010_11_001;
B[20] = 19'b00000000000_000_00_000;
B[52] = 19'b00000000000_000_00_000;
B[84] = 19'b00000000000_000_00_000;
B[116] = 19'b00000000000_000_00_000;
B[148] = 19'b01101001000_000_00_000;
B[180] = 19'b00001001000_100_00_001;
B[212] = 19'b00000000000_000_00_000;
B[244] = 19'b00000000000_000_00_000;
B[21] = 19'b00001000001_010_00_001;
B[53] = 19'b00001000011_010_00_001;
B[85] = 19'b00001000101_010_00_001;
B[117] = 19'b00001000111_010_00_001;
B[149] = 19'b00101001001_000_00_000;
B[181] = 19'b00001001001_010_00_001;
B[213] = 19'b00001001101_000_00_001;
B[245] = 19'b00001001111_010_00_001;
B[22] = 19'b00010001000_000_00_001;
B[54] = 19'b00010011000_000_00_001;
B[86] = 19'b00010101000_000_00_001;
B[118] = 19'b00010111000_000_00_001;
B[150] = 19'b10101001000_000_10_000;
B[182] = 19'b00001001000_001_10_001;
B[214] = 19'b00011101000_000_00_001;
B[246] = 19'b00011111000_000_00_001;
B[23] = 19'b00010000001_010_00_001;
B[55] = 19'b00010010011_010_00_001;
B[87] = 19'b00010100101_010_00_001;
B[119] = 19'b00010110111_010_00_001;
B[151] = 19'b11101001001_000_10_000;
B[183] = 19'b00001001001_011_10_001;
B[215] = 19'b00011101101_000_00_001;
B[247] = 19'b00011111111_010_00_001;
B[24] = 19'b00000000000_000_10_101;
B[56] = 19'b00000000000_000_10_101;
B[88] = 19'b00000000000_000_10_110;
B[120] = 19'b00000000000_000_10_110;
B[152] = 19'b01101001000_010_10_001;
B[184] = 19'b00111001000_000_10_011;
B[216] = 19'b00000000000_000_10_111;
B[248] = 19'b00000000000_000_10_111;
B[25] = 19'b00001000001_010_10_001;
B[57] = 19'b00001000011_010_10_001;
B[89] = 19'b00001000101_010_10_001;
B[121] = 19'b00001000111_010_10_001;
B[153] = 19'b00101001001_000_10_000;
B[185] = 19'b00001001001_010_10_001;
B[217] = 19'b00001001101_000_10_001;
B[249] = 19'b00001001111_010_10_001;
B[26] = 19'b00010001000_000_10_001;
B[58] = 19'b00010011000_000_10_001;
B[90] = 19'b00010101000_000_10_001;
B[122] = 19'b00010111000_000_10_001;
B[154] = 19'b10101001000_000_10_000;
B[186] = 19'b00111001000_001_10_001;
B[218] = 19'b00011101000_000_10_001;
B[250] = 19'b00011111000_000_10_001;
B[27] = 19'b00010000001_010_10_001;
B[59] = 19'b00010010011_010_10_001;
B[91] = 19'b00010100101_010_10_001;
B[123] = 19'b00010110111_010_10_001;
B[155] = 19'b11101001001_000_10_000;
B[187] = 19'b00001001001_000_10_000;
B[219] = 19'b00011101101_000_10_001;
B[251] = 19'b00011111111_010_10_001;
B[28] = 19'b00000000000_000_00_000;
B[60] = 19'b00000000000_000_00_000;
B[92] = 19'b00000000000_000_00_000;
B[124] = 19'b00000000000_000_00_000;
B[156] = 19'b01101001000_000_00_000;
B[188] = 19'b00001001000_100_00_001;
B[220] = 19'b00000000000_000_00_000;
B[252] = 19'b00000000000_000_00_000;
B[29] = 19'b00001000001_010_00_001;
B[61] = 19'b00001000011_010_00_001;
B[93] = 19'b00001000101_010_00_001;
B[125] = 19'b00001000111_010_00_001;
B[157] = 19'b00101001001_000_00_000;
B[189] = 19'b00001001001_010_00_001;
B[221] = 19'b00001001101_000_00_001;
B[253] = 19'b00001001111_010_00_001;
B[30] = 19'b00010001000_000_00_001;
B[62] = 19'b00010011000_000_00_001;
B[94] = 19'b00010101000_000_00_001;
B[126] = 19'b00010111000_000_00_001;
B[158] = 19'b10101001000_000_10_000;
B[190] = 19'b00001001000_001_10_001;
B[222] = 19'b00011101000_000_00_001;
B[254] = 19'b00011111000_000_00_001;
B[31] = 19'b00010000001_010_00_001;
B[63] = 19'b00010010011_010_00_001;
B[95] = 19'b00010100101_010_00_001;
B[127] = 19'b00010110111_010_00_001;
B[159] = 19'b11101001001_000_10_000;
B[191] = 19'b00001001001_011_10_001;
B[223] = 19'b00011101101_000_00_001;
B[255] = 19'b00011111111_010_00_001;
  end  
  wire [14:0] R = A[M[4:0]];
  reg [18:0] AluFlags;
  always @(posedge clk) if (reset) begin
    AluFlags <= 0;
  end else if (ce) begin  
    AluFlags <= B[IR];
  end

  assign Mout = {AluFlags,// 19
                 M[8:7],  // NextState // 2
                 R[14:13],// LoadT     // 2
                 R[12],   // FlagCtrl  // 1
                 R[11:7], // AddrCtrl  // 5
                 R[6:4],  // MemWrite  // 3
                 M[6:5],  // AddrBus   // 2
                 R[3:2],  // LoadPC    // 2
                 R[1:0]   // LoadSP    // 2
                 };
endmodule

