package Games;

typedef enum {MARIO, DONKEY_KONG, PACMAN, GALAGA, DEFENDER2, GOLF, PINBALL, TENNIS, EMS} game_name;

endpackage : Games